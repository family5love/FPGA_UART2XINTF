library verilog;
use verilog.vl_types.all;
entity tb_xintf_top is
end tb_xintf_top;
