library verilog;
use verilog.vl_types.all;
entity tb_xintf is
end tb_xintf;
