library verilog;
use verilog.vl_types.all;
entity tb_exe_pulse_lighting is
end tb_exe_pulse_lighting;
